module Tx(
    
);
    
endmodule